Subtrator_inst : Subtrator PORT MAP (
		clock	 => clock_sig,
		dataa	 => dataa_sig,
		datab	 => datab_sig,
		result	 => result_sig
	);
